package test_pkg;


//import uvm_pkg.sv
        import uvm_pkg::*;
//include uvm_macros.sv
        `include "uvm_macros.svh"
//`include "tb_defs.sv"
`include "source_xtn.sv"
`include "source_agent_config.sv"
`include "destination_agent_config.sv"
`include "env_config.sv"
`include "source_driver.sv"
`include "source_monitor.sv"
`include "source_sequencer.sv"
`include "source_agent.sv"
`include "source_agent_top.sv"
`include "sbase_sequence.sv"

`include "destination_xtn.sv"
`include "destination_monitor.sv"
`include "destination_sequencer.sv"
//`include "destination_sequence.sv"
`include "destination_driver.sv"
`include "destination_agent.sv"
`include "destination_agent_top.sv"
`include "dbase_sequence.sv"

`include "virtual_sequencer.sv"
`include "virtual_sequence.sv"
`include "scoreboard.sv"

`include "tb.sv"


`include "vtest_lib.sv"
endpackage
